module multiply(input logic [7:0]a, [3:0]b, output logic [7:0]c);

assign c = b*b;
endmodule

