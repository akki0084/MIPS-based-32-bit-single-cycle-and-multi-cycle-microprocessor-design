module tb();
logic clk;
logic reset;
logic [31:0] writedata;
logic [31:0]adr;
logic memwrite;
// instantiate device to be tested
TOP_M dut (clk, reset, writedata, adr, memwrite);
// initialize test
initial
begin
reset <= 1; #10; reset <= 0;
end
// generate clock to sequence tests
always
begin
clk <= 1; # 5; clk <= 0; # 5;
end
// check results
always @(negedge clk)
begin
if(memwrite) begin
if(adr===84) begin
$display ("simulation succeeded");
$stop;

end else 
if(adr!==80) begin
$display ("simulation failed");
$stop;
end
end
end
endmodule 
