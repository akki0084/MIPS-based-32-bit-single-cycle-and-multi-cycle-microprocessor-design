module CA2(input logic [7:0]A, [3:0]B, output logic [7:0]Y);
always_comb
begin
 Y[0] = A[1]? (A[0]? B[3] : B[2]) 
	    : (A[0]? B[1] : B[0]);
 Y[1] = A[2]? (A[1]? B[3] : B[2])
            : (A[1]? B[1] : B[0]);
 Y[2] = A[3]? (A[2]? B[3] : B[2])
            : (A[2]? B[1] : B[0]);
 Y[3] = A[4]? (A[3]? B[3] : B[2])
            : (A[3]? B[1] : B[0]);
 Y[4] = A[5]? (A[4]? B[3] : B[2])
            : (A[4]? B[1] : B[0]);
 Y[5] = A[6]? (A[5]? B[3] : B[2])
            : (A[5]? B[1] : B[0]);
 Y[6] = A[7]? (A[6]? B[3] : B[2])
            : (A[6]? B[1] : B[0]);
 Y[7] = A[0]? (A[7]? B[3] : B[2])
            : (A[7]? B[1] : B[0]);
end
endmodule 
